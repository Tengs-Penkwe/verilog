module my_design;
	initial begin 
		$display("Hallo Welt!");
		$finish;
	end
endmodule

